��/ / A s s e r t i o n s    
  
 / / [ 1 ]   W h e n   T e r m i n a l   C o u n t   i s   r e a c h e d   i . e .   i t   i s   a s s e r t e d   E O P n ( a c t i v e   l o w )   i s   a s s e r t e d .  
 p r o p e r t y   T e r m i n a l C o u n t _ p ;  
 d i s a b l e   i f f   ( r s t ) ;  
   @ ( p o s e d g e   c l k )  
   T C | - > ( ! E O P n )  
   e n d p r o p e r t y  
    
   T e r m i a l C o u n t _ a : a s s e r t   p r o p e r t y   T e r m i n a l C o u n t _ p ;  
    
    
    
 / / [ 2 ]   I n   s t a t e   A c t i v e   1   i f   T e r m i n a l   C o u n t   i s   r e a c h e d   N e x t   S t a t e   g o e s   t o   I n a c t i v e   0  
 p r o p e r t y   a c t i v e 1 T C _ p ;  
 d i s a b l e   i f f   ( r s t ) ;  
   @ ( p o s e d g e   c l k )  
   T C   & & ( S t a t e = = A c t i v e 1 ) | - > ( N e x t S t a t e = I n a c t i v e 0 ) ;  
   e n d p r o p e r t y  
    
   a c t i v e 1 T C _ a : a s s e r t   p r o p e r t y   a c t i v e 1 T C _ p ;  
    
    
    
 / / [ 3 ]   I n   s t a t e   A c t i v e   1   i f   T e r m i n a l   C o u n t   i s   r e a c h e d   N e x t   S t a t e   g o e s   t o   I n a c t i v e   0  
 p r o p e r t y   a c t i v e 1 T C _ p ;  
 d i s a b l e   i f f   ( r s t )  
   @ ( p o s e d g e   c l k )  
   T C   & &   ( S t a t e = = A c t i v e 1 ) | - > ( N e x t S t a t e = I n a c t i v e 0 ) ;  
   e n d p r o p e r t y  
    
   a c t i v e 1 T C _ a : a s s e r t   p r o p e r t y   a c t i v e 1 T C _ p ;  
    
    
    
 / / [ 4 ]   I n   s t a t e   A c t i v e   2   i f   T e r m i n a l   C o u n t   i s   r e a c h e d   N e x t   S t a t e   g o e s   t o   I n a c t i v e   0  
 p r o p e r t y   a c t i v e 2 T C _ p ;  
 d i s a b l e   i f f   ( r s t ) ;  
   @ ( p o s e d g e   c l k )  
   T C   & & ( S t a t e = = A c t i v e 2 ) | - > ( N e x t S t a t e = I n a c t i v e 0 ) ;  
   e n d p r o p e r t y  
    
   a c t i v e 2 T C _ a : a s s e r t   p r o p e r t y   a c t i v e 2 T C _ p ;  
    
    
    
 / / [ 5 ]   I n   s t a t e   A c t i v e   4   i f   T e r m i n a l   C o u n t   i s   r e a c h e d   N e x t   S t a t e   g o e s   t o   I n a c t i v e   0  
 p r o p e r t y   a c t i v e 2 T C _ p ;  
 d i s a b l e   i f f   ( r s t ) ;  
   @ ( p o s e d g e   c l k )  
   T C   & & ( S t a t e = = A c t i v e 4 ) | - > ( N e x t S t a t e = I n a c t i v e 0 ) ;  
   e n d p r o p e r t y  
  
   a c t i v e 4 T C _ a : a s s e r t   p r o p e r t y   a c t i v e 4 T C _ p ;  
    
    
    
 / / [ 6 ] I f   S t a t e   i s   I n a c t i v e   0   t h e n   H R Q   s h o u l d   b e   a s s e r t e d   a n d   A E N   s h o u l d   b e   d e a s s e r t e d  
 p r o p e r t y   o u t p u t I n a c t i v e 0 _ p ;  
 d i s a b l e   i f f   ( r s t )  
   @ ( p o s e d g e   c l k )  
   ( S t a t e = = I n a c t i v e 0 ) | - > ( H R Q )   & &   ( ! A E N ) ;  
   e n d p r o p e r t y  
    
   o u t p u t I n a c t i v e 0 _ a :   a s s e r t   p r o p e r t y   o u t p u t I n a c t i v e 0 _ p ;  
    
    
    
 / / [ 7 ] I f   s t a t e   i s   A c t i v e   1   t h e n   A E N   A D S T B   l d U p p e r A d d r   D A C K   s h o u l d   b e   a s s e r t e d  
 p r o p e r t y   o u t p u t A c t i v e 1 _ p ;  
 d i s a b l e   i f f ( r s t )  
 @ ( p o s e d g e   c l k )  
 ( S t a t e = = A c t i v e 1 ) | = > ( A E N )   & &   ( A D S T B )   & &   ( l d U p p e r A d d r e s s )   & &   ( D A C K ) ;  
 e n d p r o p e r t y  
  
 o u t p u t A c t i v e 1 _ a : a s s e r t   p r o p e r t y   o u t p u t A c t i v e 1 _ p ;  
  
  
  
 / / [ 8 ] I f   s t a t e   i s   A c t i v e   2   t h e n   A D S T B   a n d   l d U p p e r A d d r   s h o u l d   b e   d e a s s e r t e d  
 p r o p e r t y   o u t p u t A c t i v e 2 _ p ;  
 d i s a b l e   i f f ( r s t )  
 @ ( p o s e d g e   c l k )  
 ( S t a t e = = A c t i v e 2 ) | - > ( A D S T B )   & &   ( ! l d U p p e r A d d r e s s )  
 e n d p r o p e r t y  
  
 o u t p u t A c t i v e 2 _ a : a s s e r t   p r o p e r t y   o u t p u t A c t i v e 2 _ p ;  
  
  
  
 / / [ 9 ] I f   s t a t e   i s   I n a c t i v e 0   t h e n   c h e c k   N e x t   S t a t e  
 p r o p e r t y   n e x t s t a t e I n a c t i v e 0 _ p ;  
 d i s a b l e   i f f ( r s t )  
 @ ( p o s e d g e   c l k )  
 c h i p S e l N   & &   D R E Q   & &   ( S t a t e = I n a c t i v e 0 ) | = > ( N e x t S t a t e = A c t i v e 0 ) ;  
 e n d p r o p e r t y  
  
 n e x t s t a t e I n a c t i v e 0 _ a :   a s s e r t   p r o p e r t y   n e x t s t a t e I n a c t i v e 0 _ p ;  
  
  
  
 / / [ 1 0 ] I f   s t a t e   i s   A c t i v e   0   t h e n   c h e c k   N e x t   S t a t e  
 p r o p e r t y   n e x t s t a t e A c t i v e 0 _ p ;  
 d i s a b l e   i f f ( r s t )  
 @ ( p o s e d g e   c l k )  
 H L D A   & &   ( S t a t e = A c t i v e 0 ) | = > ( N e x t S t a t e = A c t i v e 1 ) ;  
 e n d p r o p e r t y  
  
 n e x t s t a t e A c t i v e 0 _ a :   a s s e r t   p r o p e r t y   n e x t s t a t e A c t i v e 0 _ p ;  
  
  
  
 / / [ 1 1 ] I f   s t a t e   i s   A c t i v e   1   t h e n   c h e c k   N e x t   S t a t e  
 p r o p e r t y   n e x t s t a t e A c t i v e 1 _ p ;  
 d i s a b l e   i f f ( r s t )  
 @ ( p o s e d g e   c l k )  
 E O P n   & &   ( S t a t e = A c t i v e 1 )   | = > ( N e x t S t a t e = A c t i v e 2 ) ;  
 e n d p r o p e r t y  
  
 n e x t s t a t e A c t i v e 1 _ a :   a s s e r t   p r o p e r t y   n e x t s t a t e A c t i v e 1 _ p ;  
  
  
  
 / / [ 1 2 ] I f   s t a t e   i s   A c t i v e   2   t h e n   c h e c k   N e x t   S t a t e    
 p r o p e r t y   n e x t s t a t e A c t i v e 4 _ p ;  
 d i s a b l e   i f f ( r s t )  
 @ ( p o s e d g e   c l k )  
 E O P n   & &   ( S t a t e = A c t i v e 2 ) | = > ( N e x t S a t e = A c t i v e 4 ) ;  
 e n d p r o p e r t y  
  
 n e x t s t a t e A c t i v e 2 _ a :   a s s e r t   p r o p e r t y   n e x t s t a t e A c t i v e 2 _ p ;  
  
  
  
 / / [ 1 3 ] I f   s t a t e   i s   A c t i v e   4   t h e n   c h e c k   N e x t   S t a t e   i f   c a r r y   p r e s e n t  
 p r o p e r t y   c a r r y P r e s e n t A c t i v e 4 _ p ;  
 d i s a b l e   i f f ( r s t )  
 @ ( p o s e d g e   c l k )  
 c a r r y P r e s e n t   & &   ( S t a t e = A c t i v e 4 ) | = > ( N e x t S a t e = A c t i v e 1 ) ;  
 e n d p r o p e r t y  
  
 c a r r y P r e s e n t A c t i v e 4 _ a :   a s s e r t   p r o p e r t y   c a r r y P r e s e n t A c t i v e 4 _ p ;  
  
  
  
 / / [ 1 4 ] I f   s t a t e   i s   A c t i v e   4   t h e n   c h e c k   N e x t   S t a t e   i f   n o   c a r r y   p r e s e n t    
 p r o p e r t y   n o C a r r y A c t i v e 4 _ p ;  
 d i s a b l e   i f f ( r s t )  
 @ ( p o s e d g e   c l k )  
 ( ! c a r r y P r e s e n t )   & &   ( S t a t e = A c t i v e 4 )   | = > ( N e x t S t a t e = A c t i v e 2 ) ;  
 e n d p r o p e r t y  
  
 n o C a r r y A c t i v e 4 _ a :   a s s e r t   p r o p e r t y   n o C a r r y A c t i v e 4 _ p ;  
  
  
  
 / / [ 1 5 ] I f   A d d r e s s   S t r o b e   i s   h i g h   f o r   o n l y   o n e   c y c l e  
  
 p r o p e r t y   A d d r e s s S t r o b e _ p ;  
 d i s a b l e   i f f ( r s t )  
 	 @ ( p o s e d g e   c l k )  
 	 c h i p S e l N   | - >   A D S T B   # # 1   ( ~ A D S T B ) ;  
 e n d p r o p e r t y  
  
 A d d r e s s S t r o b e _ a :   a s s e r t   p r o p e r t y   ( A d d r e s s S t r o b e _ p ) ;  
  
  
  
 / / [ 1 6 ]   E O P n   i s   d e a s s e r t e d   w h e n   t r a n s f e r   i s   c o m p l e t e  
  
 p r o p e r t y   E O P C h e c k _ p ;  
 d i s a b l e   i f f ( r s t )  
 	 @ ( p o s e d g e   c l k )  
 	 ( ( c h i p S e l N )   & &   ( T C ) )   | = >   ( ! E O P n ) ;  
 e n d p r o p e r t y  
  
 E O P C h e c k _ a :   a s s e r t   p r o p e r t y   ( E O P C h e c k _ p ) ;  
  
  
  
 / / [ 1 7 ]     W h e n   S t a t e   i s   A c t i v e   4   a n d   i s R e a d   i s   z e r o   t h e n   M E M W n   a n d   I O R n   a r e   a s s e r t e d   ( a c t i v e   l o w )  
 p r o p e r t y   i s R e a d z e r o _ p ;  
 d i s a b l e   i f f ( r s t )  
 	 @ ( p o s e d g e   c l k )  
 	     ( S t a t e = = A c t i v e 4 )   & &   ( i s R e a d = = 0 ) | - > ( ! M E M W n )   & &   ( ! I O R n )  
 e n d p r o p e r t y  
  
 i s R e a d z e r o _ a :   a s s e r t   p r o p e r t y   ( i s R e a d z e r o _ p ) ;  
  
  
  
 / / [ 1 8 ]     W h e n   S t a t e   i s   A c t i v e   4   a n d   i s R e a d   i s   o n e   t h e n   M E M R n   a n d   I O W n   a r e   a s s e r t e d   ( a c t i v e   l o w )  
 p r o p e r t y   i s R e a d o n e _ p ;  
 d i s a b l e   i f f ( r s t )  
 	 @ ( p o s e d g e   c l k )  
 	     ( S t a t e = = A c t i v e 4 )   & &   ( i s R e a d = = 1 ) | - > ( ! M E M R n )   & &   ( ! I O W n )  
 e n d p r o p e r t y  
  
 i s R e a d o n e _ a :   a s s e r t   p r o p e r t y   ( i s R e a d o n e _ p ) ;  
  
  
  
  
  
    
   